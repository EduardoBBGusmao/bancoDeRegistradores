module readregister(Q, );