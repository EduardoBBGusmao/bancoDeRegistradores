module reg_zero(Q);
 output wire [31:0] Q;
 assign Q = 32'b0;
endmodule